Temporary first version.
